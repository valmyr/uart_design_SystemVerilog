module


parameterizedCounter(.pMODULE(pMODULE),.WIDTH(WIDTH))overSamplingCounter(
    .nreset(nreset),
    .clock (clock),
    .start (start1_counter),
    .done  (done1_counter)
);


endmodule